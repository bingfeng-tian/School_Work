module dec_7seg (D, Q1, Q2);
input   [3:0]D;
output  [6:0]Q1, Q2;
reg     [6:0]Q1, Q2;

always@(D)
    if      (D==4'b0000)    Q1 = 7'b0000001;
    else if (D==4'b0001)    Q1 = 7'b1001111;
    else if (D==4'b0010)    Q1 = 7'b0010010;
    else if (D==4'b0011)    Q1 = 7'b0000110;
    else if (D==4'b0100)    Q1 = 7'b1001100;
    else if (D==4'b0101)    Q1 = 7'b0100100;
    else if (D==4'b0110)    Q1 = 7'b0100000;
    else if (D==4'b0111)    Q1 = 7'b0001101;
    else if (D==4'b1000)    Q1 = 7'b0000000;
    else if (D==4'b1001)    Q1 = 7'b0000100;
    else if (D==4'b1010)    Q1 = 7'b0001000;
    else if (D==4'b1011)    Q1 = 7'b1100000;
    else if (D==4'b1100)    Q1 = 7'b0110001;
    else if (D==4'b1101)    Q1 = 7'b1000010;
    else if (D==4'b1110)    Q1 = 7'b0110000;
    else                    Q1 = 7'b0111000;

always@(D)
    case(D)
        (4'b0000):      Q2 = 7'b0000001;
        (4'b0001):      Q2 = 7'b1001111;
        (4'b0010):      Q2 = 7'b0010010;
        (4'b0011):      Q2 = 7'b0000110;
        (4'b0100):      Q2 = 7'b1001100;
        (4'b0101):      Q2 = 7'b0100100;
        (4'b0110):      Q2 = 7'b0100000;
        (4'b0111):      Q2 = 7'b0001101;
        (4'b1000):      Q2 = 7'b0000000;
        (4'b1001):      Q2 = 7'b0000100;
        (4'b1010):      Q2 = 7'b0001000;
        (4'b1011):      Q2 = 7'b1100000;
        (4'b1100):      Q2 = 7'b0110001;
        (4'b1101):      Q2 = 7'b1000010;
        (4'b1110):      Q2 = 7'b0110000;
        default:        Q2 = 7'b0111000;
    endcase


endmodule